* Atmega simple signal gen
* connections:      Pwr
*                   |   Gnd
*                   |   |   B0  .... B
*                   |   |   |
.SUBCKT atmega      1   2   3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
*RLoad 1 2 30
VGenB 60 0 Pulse(0 3.3 0 0.00001 0.00001 0.0001 0.0002)
VGenC 70 0 Pulse(0 3.3 0 0.00001 0.00001 0.0002 0.0004)
R0 60 3 100
R1 60 4 100
R2 60 5 100
R3 60 6 100
R4 60 7 100
R5 60 8 100
R6 60 9 100
R7 60 10 100
R10 70 11 100
R11 70 12 100
R12 70 13 100
R13 70 14 100
R14 70 15 100
R15 70 16 100
R16 70 17 100
R17 70 18 100
R19 70 19 100
R20 70 20 100
R21 70 21 100
R22 70 22 100
R23 70 23 100
R24 70 24 100
R25 70 25 100
R26 70 26 100
.ENDS atmega
