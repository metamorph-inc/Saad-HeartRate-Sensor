*************************************************************
* Ngspice .cir file for C_TANT_1210_220u_6.3V_20%_AVX
*************************************************************
* AVX Tantalum Capacitor TLJT227K006R2000
*
.SUBCKT TLJT227K006R2000 POS NEG

*PARASITIC INDUCTANCE
LESL POS 2 1.800000E-009
RELS POS 2 10

*LEAKAGE CURRENT & REVERSE BIAS EFFECTS
RP 2 NEG 5.000000E+005
DP NEG 2 DFWD

*RC-LADDER MODEL OF FREQUENCY EFFECTS
R1 2 3 RMOD1 1.899567E-001
C1 2 3 CMOD1 1.852467E-003
R2 3 4 RMOD2 2.512347E-001
C2 4 NEG CMOD2 7.171424E-006
R3 4 5 RMOD3 1.539633E-001
C3 5 NEG CMOD3 1.434285E-005
R4 5 6 RMOD4 2.282102E-001
C4 6 NEG CMOD4 2.868570E-005
R5 6 7 RMOD5 3.447706E-001
C5 7 NEG CMOD5 5.737139E-005
R6 7 8 RMOD6 6.200312E-001
C6 8 NEG CMOD6 1.147428E-004

.MODEL CMOD1 C (TNOM=25 TC1=1.463615E-003 TC2=-4.147800E-005)
.MODEL CMOD2 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL CMOD3 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL CMOD4 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL CMOD5 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL CMOD6 C (TNOM=25 TC1=3.749220E-004 TC2=2.806000E-006)
.MODEL RMOD1 R (TNOM=25 TC1=5.948893E-003 TC2=5.337100E-005)
.MODEL RMOD2 R (TNOM=25 TC1=-1.770874E-003 TC2=1.281300E-005)
.MODEL RMOD3 R (TNOM=25 TC1=-7.138201E-003 TC2=2.153200E-005)
.MODEL RMOD4 R (TNOM=25 TC1=-7.138201E-003 TC2=2.153200E-005)
.MODEL RMOD5 R (TNOM=25 TC1=-7.138201E-003 TC2=2.153200E-005)
.MODEL RMOD6 R (TNOM=25 TC1=-7.138201E-003 TC2=2.153200E-005)
.MODEL DFWD D (RS=0.1 IS=8E-7 N=2.5 XTI=0 EG=0.1)

.ENDS TLJT227K006R2000
*************************************************************
